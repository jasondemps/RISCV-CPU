library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all
--
--  package Utility
--  -- Was working on unsigned -> signed in 1 function...
--end Utility;
--
--package body Utility
--begin
--
--end Utility;
