library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

use work.declares.all;

package instr_set is

end instr_set;

package body instr_set is



end instr_set;
