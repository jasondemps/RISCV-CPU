library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.declares.all;

entity CPU is
  port(
    clock : in std_logic;
    
    );
end CPU;

architecture Sim_CPU of CPU is

begin

  -- FETCH
  process(clock)
  begin

    
    
    end process;

  

end Sim_CPU;
