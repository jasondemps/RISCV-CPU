library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Branch_Predict is
  port (

);
end Branch_Predict;

architecture Sim_Branch_Predict of Branch_Predict is

begin


end Sim_Branch_Predict;
